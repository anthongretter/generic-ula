-- arquivo que juntara BO e BC de ula, com saidas PQ, S e flagZ.