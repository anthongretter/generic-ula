-- bloco de controle ula;; enA, enB, enPC, enOut, opcode, etc.