-- contem: regpc, mem_dados, regA, regB, regOP; ula inicial, regpq, regs, regz.